module Prio_Enco(i,y,z);
input [22:0]i;
output [4:0]y;
output z;

assign z= i[0] | i[1] | i[2] | i[3] | i[4] | i[5] | i[6] | i[7] | i[8]|i[9]|i[10]|i[11]|i[12]|i[13]|i[14]|i[15] | i[16]|i[17]|i[18]|i[19]|i[20]|i[21]|i[22];
assign y[4]=i[22]|i[21]|i[20]|i[19]|i[18]|i[17]|i[16];
assign y[3]=~i[22] & ~i[21] & ~i[20] & ~i[19] & ~i[18] & ~i[17] & ~i[16]  & (i[15] | i[14] | i[13] | i[12] | i[11] | i[10] | i[9] | i[8]);
assign y[2]=i[22] | i[21] | i[20] | (~i[19] & ~i[18] & ~i[17] & ~i[16]) & (i[15] | i[14] | i[13] | i[12] | (~i[11] & ~i[10] & ~i[9] & ~i[8]) & (i[7] | i[6] | i[5] | i[4]));
assign y[1]=i[22] | (~i[21] & ~i[20]) & (i[19] | i[18]) | (~i[21] & ~i[20] & ~i[17] & ~i[16]) & (i[15] | i[14]) | (~i[21] & ~i[20] & ~i[17] & ~i[16] & ~i[13] & ~i[12]) & (i[11] | i[10]) | (~i[21] & ~i[20] & ~i[17] & ~i[16] & ~i[13] & ~i[12] & ~i[9] & ~i[8]) & ((i[7] | i[6]) | (~i[5] & ~i[4]) & (i[3] & i[2]));
assign y[0]=~i[22] & (i[21] | ~i[20] & (i[19] | ~i[18] & (i[17] | ~i[16] & (i[15] | ~i[14] & (i[13] | ~i[12] & (i[11] | ~i[10] & (i[9] | ~i[8] & (i[7] | ~i[6] & (i[5] | ~i[4] & (i[3] | ~i[2] & (i[1])))))))))));

endmodule
