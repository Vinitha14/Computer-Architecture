`include "FM.v"
module IEEEFM_tb;
reg [15:0]a; reg[15:0]b;
wire [15:0]y;
wire [32:0]y1;

initial begin
$dumpfile("IEEEFM.vcd");
$dumpvars(0,IEEEFM_tb);
$display("a      			   b			 y");
$monitor("%b,  %b, %b", a, b,y);
end

initial begin
a=16'b0100101110000000;b=16'b0100001000000000; //15,3 = 45
#20 a=16'b0100101110000000;b=16'b1100001000000000;//15,-3
#20 a=16'b1100101110000000;b=16'b0100001000000000;//-15,3
#20 a=16'b1100101110000000;b=16'b1100001000000000;//-15,-3

#20 a=16'b0100001000000000;b=16'b1100101110000000;//3,-15
#20 a=16'b0100001000000000;b=16'b0100101110000000;//3,15

#20 a=16'b0100101110000000;b=16'b0100101110000000;//15,15
#20 a=16'b0100101110000000;b=16'b1100101110000000;//15,-15
#20 a=16'b1100101110000000;b=16'b0100101110000000;//-15,15
#20 a=16'b1100101110000000;b=16'b1100101110000000;//-15,-15

#20 a=16'b0100100010000000;b=16'b0100100000000000;//9,8
#20 a=16'b0100100010000000;b=16'b1100100000000000;//9,-8
#20 a=16'b1100100010000000;b=16'b0100100000000000;//-9,8
#20 a=16'b1100100010000000;b=16'b1100100000000000;//-9,-8

#20 a=16'b0011100000000000;b=16'b0100101000100110;//0.5,12.3 = 16.5
#20 a=16'b0011100000000000;b=16'b1100101000100110;//0.5,-12.3
#20 a=16'b1011100000000000;b=16'b0100101000100110;//-0.5,12.3
#20 a=16'b1011100000000000;b=16'b1100101000100110;//-0.5,-12.3

#20 a=16'b0100101110000000;b=16'b0000000000000000;//15,0
#20 a=16'b0000000000000000;b=16'b1100101110000000;//0,-15

#20 a=16'b0000000000000000;b=16'b0000000000000000;//0,0
end

FM obj(
.a(a),
.b(b),
.y(y),
.y1(y1)
);

initial
#1000 $finish;
endmodule
