`include "floating.v"
module IEEEfloatingpt_tb;
reg [15:0]C;
reg[15:0]D;
reg ch;
wire [15:0]A;

initial begin
$dumpfile("IEEEfloating.vcd");
$dumpvars(0,IEEEfloatingpt_tb);
$display("C      		   D		    ch  A");
$monitor("%b,  %b, %b, %b", C, D,ch, A);
end

initial begin
    C=16'b0100101110000000;D=16'b0100001000000000; ch=0;//15,3
#20 C=16'b0100101110000000;D=16'b1100001000000000; ch=0; //15,-3
#20 C=16'b1100101110000000;D=16'b0100001000000000; ch=0;//-15,3
#20 C=16'b1100101110000000;D=16'b1100001000000000; ch=0;//-15,-3

#20 C=16'b0100001000000000;D=16'b1100101110000000; ch=0; //3,-15
#20 C=16'b0100001000000000;D=16'b1100101110000000; ch=1;//3,-15
#20 C=16'b0100001000000000;D=16'b0100101110000000; ch=0; //3,15
#20 C=16'b0100001000000000;D=16'b0100101110000000; ch=1;//3,15

#20 C=16'b0100101110000000;D=16'b0100001000000000; ch=1;//15,3
#20 C=16'b0100101110000000;D=16'b1100001000000000; ch=1; //15,-3
#20 C=16'b1100101110000000;D=16'b0100001000000000; ch=1;//-15,3
#20 C=16'b1100101110000000;D=16'b1100001000000000; ch=1;//-15,-3

#20 C=16'b0011100000000000;D=16'b0100101000100110; ch=1; //0.5,12.3
#20 C=16'b0011100000000000;D=16'b1100101000100110; ch=1;//0.5,-12.3
#20 C=16'b1011100000000000;D=16'b0100101000100110; ch=1;//-0.5,12.3
#20 C=16'b1011100000000000;D=16'b1100101000100110; ch=1;//-0.5,-12.3

#20 C=16'b0011100000000000;D=16'b0100101000100110; ch=0; //0.5,12.3
#20 C=16'b0011100000000000;D=16'b1100101000100110; ch=0;//0.5,-12.3
#20 C=16'b1011100000000000;D=16'b0100101000100110; ch=0;//-0.5,12.3
#20 C=16'b1011100000000000;D=16'b1100101000100110; ch=0;//-0.5,-12.3

#20 C=16'b0100101110000000;D=16'b0100101110000000; ch=0;//15,15
#20 C=16'b0100101110000000;D=16'b1100101110000000; ch=0;//15,-15
#20 C=16'b1100101110000000;D=16'b0100101110000000; ch=0;//-15,15
#20 C=16'b1100101110000000;D=16'b1100101110000000; ch=0;//-15,-15

#20 C=16'b0100101110000000;D=16'b0100101110000000; ch=1;//15,15
#20 C=16'b0100101110000000;D=16'b1100101110000000; ch=1;//15,-15
#20 C=16'b1100101110000000;D=16'b0100101110000000; ch=1;//-15,15
#20 C=16'b1100101110000000;D=16'b1100101110000000; ch=1;//-15,-15

#20 C=16'b0100100010000000;D=16'b0100100000000000; ch=0;//9,8
#20 C=16'b0100100010000000;D=16'b1100100000000000; ch=0;//9,-8
#20 C=16'b1100100010000000;D=16'b0100100000000000; ch=0;//-9,8
#20 C=16'b1100100010000000;D=16'b1100100000000000; ch=0;//-9,-8

#20 C=16'b0100100010000000;D=16'b0100100000000000; ch=1;//9,8
#20 C=16'b0100100010000000;D=16'b1100100000000000; ch=1;//9,-8
#20 C=16'b1100100010000000;D=16'b0100100000000000; ch=1;//-9,8
#20 C=16'b1100100010000000;D=16'b1100100000000000; ch=1;//-9,-8

#20 C=16'b0100101110000000;D=16'b0000000000000000; ch=0;//15,0
#20 C=16'b0000000000000000;D=16'b1100101110000000; ch=0;//0,-15
#20 C=16'b0100101110000000;D=16'b0000000000000000; ch=1;//15,0
#20 C=16'b0000000000000000;D=16'b1100101110000000; ch=1;//0,-15

#20 C=16'b0000000000000000;D=16'b0000000000000000; ch=0;//0,0
#20 C=16'b0000000000000000;D=16'b0000000000000000; ch=1;//0,0

end

IEEEfloatingpt addsub(
.C(C),
.D(D),
.ch(ch),
.A(A)
);

initial
#1000 $finish;
endmodule
